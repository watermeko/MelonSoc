parameter M=32;
parameter N=32;
parameter MSB=32;
parameter LATENCY=2;
